//module base (input [2:0] rng,
//				  input [9:0] blockX, blockY, blockS,
//					output [9:0] shapeX, shapeY, shapeS);
//					
//			
//
//always_comb
//	begin
//		unique case (rng)
//		// I
//		3'b000 : 
//		// J
//		3'b001 : 
//		// L
//		3'b010 :
//		// S
//		3'b100 :
//		// Z
//		3'b011 :
//		// T
//		3'b110 :
//		// O
//		3'b111 :
//		
//	end
//	
//	
//endmodule
//
//module rotations (input [7:0] keycode, input [2:0] rng, 
//						output [9:0] shapeX, shapeY, shapeS);
//
//
//// predraw rotations
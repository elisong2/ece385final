module block (input frameClk, reset, 
				  output [9:0] blockX, blockY);
				  
				  
endmodule